`define FV_RIDECORE_INSERT_FV
`define FV_SUPER_SCALAR_2 
