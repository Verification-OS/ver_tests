`define FV_DUT_INSERT_FV

`define RV32E 0
`define RV32M 1

`define FV_TRIM_INDIVIDUAL_INSTRUCTIONS_CVA6
