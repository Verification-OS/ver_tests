`define FV_DUT_INSERT_FV

`define NR_LANES 4
`define RVV_ARIANE 1'b1
`define VLEN (`NR_LANES*8*64)

`define RV32E 0
`define RV32M 1

`define FV_TRIM_INDIVIDUAL_INSTRUCTIONS_4
