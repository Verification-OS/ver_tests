// use the same define for insertion in riscy nd zeroriscy to keep the RTL code more similar
`define FV_RISCY_INSERT_FV
// define that selects the core in riscy_wrapper (shared b.w. zeroriscy and riscy)
`define USE_FOR_RISCY

`define RV32E 0
`define RV32M 1

`define FV_TRIM_INDIVIDUAL_INSTRUCTIONS_4
